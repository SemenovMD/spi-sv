package axil_pkg;

    parameter                               AXI_DATA_WIDTH                  = 32;
    parameter                               AXI_ADDR_WIDTH                  = 32;

    parameter                               CLOCK                           = 100_000_000;
    parameter                               SPI_FREQ                        = 5_000_000;

endpackage
